module two(inputA, shift_clk, latch_clk, reset, output_enable, SQ, QA, QB, QC, QD, QE, QF, QG, QH);
input inputA, shift_clk, latch_clk, reset, output_enable;
output SQ, QA, QB, QC, QD, QE, QF, QG, QH;

//your code~~

endmodule